module top(output q);
assign q = 1'b1;
endmodule
