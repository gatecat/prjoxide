
(* \db:architecture ="LFCPNX", \db:device ="LFCPNX-100", \db:package ="LFG672", \db:speed ="7_High-Performance_1.0V", \db:timestamp =1576073342, \db:view ="physical" *)
module top (
    
);
    (* \dm:cellmodel_primitives ="K0=i48_3_lut", \dm:primitive ="SLICE", \dm:programming ="MODE:${mode} ${config}", \dm:site ="R2C2${z}" *) 
    SLICE SLICE_I ( );
endmodule
